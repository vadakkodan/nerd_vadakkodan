library verilog;
use verilog.vl_types.all;
entity siso_book_tb is
end siso_book_tb;
